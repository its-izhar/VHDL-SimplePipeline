-- Greg Stitt
-- University of Florida

library ieee;
use ieee.std_logic_1164.all;

use work.config_pkg.all;
use work.user_pkg.all;

entity user_app is
    port (
        clk : in std_logic;
        rst : in std_logic;

        -- memory-map interface
        mmap_wr_en   : in  std_logic;
        mmap_wr_addr : in  std_logic_vector(MMAP_ADDR_RANGE);
        mmap_wr_data : in  std_logic_vector(MMAP_DATA_RANGE);
        mmap_rd_en   : in  std_logic;
        mmap_rd_addr : in  std_logic_vector(MMAP_ADDR_RANGE);
        mmap_rd_data : out std_logic_vector(MMAP_DATA_RANGE)
        );
end user_app;

architecture default of user_app is

    signal go   : std_logic;
    signal size : std_logic_vector(C_MEM_ADDR_WIDTH downto 0);
    signal done : std_logic;

    signal mem_in_wr_data       : std_logic_vector(C_MEM_IN_WIDTH-1 downto 0);
    signal mem_in_wr_addr       : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal mem_in_rd_data       : std_logic_vector(C_MEM_IN_WIDTH-1 downto 0);
    signal mem_in_rd_addr       : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal mem_in_wr_en         : std_logic;
    signal mem_in_rd_addr_valid : std_logic;

    signal mem_out_wr_data       : std_logic_vector(C_MEM_OUT_WIDTH-1 downto 0);
    signal mem_out_wr_addr       : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal mem_out_rd_data       : std_logic_vector(C_MEM_OUT_WIDTH-1 downto 0);
    signal mem_out_rd_addr       : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal mem_out_wr_en         : std_logic;
    signal mem_out_wr_data_valid : std_logic;
    signal mem_out_done          : std_logic;
    
    --I/P Addr generator
    signal ip_addr_gen_rd_addr   : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal ip_addr_gen_valid_out, ip_addr_gen_sel_mux_in   : std_logic;
    
    --Pipeline
    signal pipeline_valid_out   : std_logic;
    signal pipeline_data_out    : std_logic_vector(C_MEM_OUT_WIDTH-1 downto 0);

    --O/P Addr generator
    signal op_addr_gen_wr_addr   : std_logic_vector(C_MEM_ADDR_WIDTH-1 downto 0);
    signal op_addr_gen_wr_en   : std_logic;
    
	signal ip_addr_gen_mode_out 	: std_logic;     -- 0: Read Mode, 1: Write Mode
    signal op_addr_gen_mode_out    : std_logic;
    
    signal ip_addr_gen_size_out     : std_logic_vector(C_MEM_ADDR_WIDTH downto 0);
    signal op_addr_gen_size_out     : std_logic_vector(C_MEM_ADDR_WIDTH downto 0);   

    signal ip_addr_gen_go        : std_logic;
    signal op_addr_gen_go        : std_logic;

    signal ip_addr_gen_done    : std_logic    := '0';
    signal op_addr_gen_done    : std_logic    := '0';   

	-- Muxes
	signal mux1_out : std_logic_vector(C_MEM_IN_WIDTH downto 0) := (others => '0');
	signal mux2_out : std_logic_vector(C_MEM_OUT_WIDTH downto 0) := (others => '0');

begin

	------------------------------------------------------------------------------
    U_MMAP : entity work.memory_map
        port map (
            clk     => clk,
            rst     => rst,
            wr_en   => mmap_wr_en,
            wr_addr => mmap_wr_addr,
            wr_data => mmap_wr_data,
            rd_en   => mmap_rd_en,
            rd_addr => mmap_rd_addr,
            rd_data => mmap_rd_data,
		
			-- TODO: connect to appropriate logic
            go              => go,         
            size            => size,       
            done            => done,       
			
			-- already connected to block RAMs
			-- the memory map functionality writes to the input ram
			-- and reads from the output ram
            mem_in_wr_data  => mem_in_wr_data,
            mem_in_wr_addr  => mem_in_wr_addr,
            mem_in_wr_en    => mem_in_wr_en,
            mem_out_rd_data => mem_out_rd_data,
            mem_out_rd_addr => mem_out_rd_addr
            );
	------------------------------------------------------------------------------

	U_CONTROLLER : entity work.controller
		port map (
			clk	=> clk,
			rst => rst,
       
			-- Mode control out for address generators
            ip_addr_gen_mode_out => ip_addr_gen_mode_out,
            op_addr_gen_mode_out => op_addr_gen_mode_out,

            -- Size of memory (i.e. The number of addressess to be generated by Address Generator)
            ip_addr_gen_size_out => ip_addr_gen_size_out,
            op_addr_gen_size_out => op_addr_gen_size_out,
               
            -- Address Generators Control I/O
            ip_addr_gen_go => ip_addr_gen_go,
            op_addr_gen_go => op_addr_gen_go,
            ip_addr_gen_done => ip_addr_gen_done,
            op_addr_gen_done => op_addr_gen_done,

			-- Controller Control I/O
			go => go,
			done => done,

			-- Size in for controller
			size => size );

	------------------------------------------------------------------------------
    -- input address generator (READ Mode)
    -- read from input memory
    -- data out to datapath from input memory
    U_ADDR_GEN_IN : entity work.addr_generator(default)
        generic map (
            ADDR_WIDTH  => C_MEM_ADDR_WIDTH)
        port map (
            clk   => clk,
            rst   => rst,
            start => ip_addr_gen_go, --from controller //DONE
            done  => ip_addr_gen_done, --to controller //DONE
            mode  => ip_addr_gen_mode_out,       -- READ Mode, from controller //DONE
            size  => ip_addr_gen_size_out,       -- from controller //DONE
			pipeIn_mux_sel => ip_addr_gen_sel_mux_in,
            valid_in => '0',
            valid_out => ip_addr_gen_valid_out,
            rd_addr  => ip_addr_gen_rd_addr);
	------------------------------------------------------------------------------

	
	------------------------------------------------------------------------------
    -- input memory
    -- written to by memory map
    -- read from by controller+datapath
    U_MEM_IN : entity work.ram(SYNC_READ)
        generic map (
            num_words  => 2**C_MEM_ADDR_WIDTH,
            word_width => C_MEM_IN_WIDTH,
            addr_width => C_MEM_ADDR_WIDTH)
        port map (
            clk   => clk,
            wen   => mem_in_wr_en,
            waddr => mem_in_wr_addr,
            wdata => mem_in_wr_data,
            raddr => ip_addr_gen_rd_addr,  -- TODO: connect to input address generator //DONE
            rdata => mem_in_rd_data); -- TODO: connect to pipeline input //DONE
	------------------------------------------------------------------------------

	------------------------------------------------------------------------------
    -- input mux to pipeline (Muxes data and valid_out together)
    -- input from data read from input memory
    -- output to datapath
	-- select is controlled from input address generator
	U_MUX_IN : entity work.mux_2x1(WITH_SELECT)
		generic map( DATA_WIDTH => C_MEM_IN_WIDTH )
		port map (
			in1 => (others => '0'),
			in2(C_MEM_IN_WIDTH-1 downto 0) => mem_in_rd_data(C_MEM_IN_WIDTH-1 downto 0),
			in2(C_MEM_IN_WIDTH) => ip_addr_gen_valid_out,
			sel => ip_addr_gen_sel_mux_in,
			output(C_MEM_IN_WIDTH-1 downto 0) => mux1_out(C_MEM_IN_WIDTH-1 downto 0),
			output(C_MEM_IN_WIDTH) => mux1_out(C_MEM_IN_WIDTH)
		);	
	------------------------------------------------------------------------------
	
	------------------------------------------------------------------------------
    -- PIPELINE
    -- data from input memory
    -- data out to output memory
    U_PIPELINE : entity work.datapath(default)
        generic map (
            data_width_in  => C_MEM_IN_WIDTH,
            data_width_out => C_MEM_OUT_WIDTH )
        port map (
            pipe_clk   => clk,
            pipe_rst   => rst,
            pipe_en    => '1',
            valid_in(0)   => mux1_out(C_MEM_IN_WIDTH),			-- from mux (MSB)
            valid_out(0) => pipeline_valid_out,
            pipe_data_in    => mux1_out(C_MEM_IN_WIDTH-1 downto 0),		-- from mux (MSB-1....0)
            pipe_data_out   => pipeline_data_out);
	------------------------------------------------------------------------------

	------------------------------------------------------------------------------
    -- output mux at pipeline output (Muxes data and valid_out together)
    -- input from pipeline
    -- output to output memory	
	-- select is controlled by write enable from output address generator
	U_MUX_OUT : entity work.mux_2x1(WITH_SELECT)
		generic map( DATA_WIDTH => C_MEM_OUT_WIDTH )
		port map (
			in1 => (others => '0'),
			in2(C_MEM_OUT_WIDTH-1 downto 0) => pipeline_data_out,
			in2(C_MEM_OUT_WIDTH) => pipeline_valid_out,
			sel => op_addr_gen_wr_en,									-- wr_en from output addr_generator
			output(C_MEM_OUT_WIDTH-1 downto 0) => mux2_out(C_MEM_OUT_WIDTH-1 downto 0),
			output(C_MEM_OUT_WIDTH) => mux2_out(C_MEM_OUT_WIDTH)
		);	
	------------------------------------------------------------------------------
	
	------------------------------------------------------------------------------
    -- output address generator (WRITE Mode)
    -- write to output memory
    -- data in from datapath to output memory
    U_ADDR_GEN_OUT : entity work.addr_generator(default)
        generic map (
            ADDR_WIDTH  => C_MEM_ADDR_WIDTH)
        port map (
            clk   => clk,
            rst   => rst,
            start => op_addr_gen_go, --from controller //DONE
            done  => op_addr_gen_done, --to controller //DONE
            mode  => op_addr_gen_mode_out,      -- WRITE Mode, from Controller //DONE
            size  => op_addr_gen_size_out,      -- from controller //DONE
            valid_in => pipeline_valid_out,
            wr_en   => op_addr_gen_wr_en,
            wr_addr  => op_addr_gen_wr_addr ); 
	------------------------------------------------------------------------------

	
	------------------------------------------------------------------------------
    -- output memory
    -- written to by controller+datapath
    -- read from by memory map
    U_MEM_OUT : entity work.ram(SYNC_READ)
        generic map (
            num_words  => 2**C_MEM_ADDR_WIDTH,
            word_width => C_MEM_OUT_WIDTH,
            addr_width => C_MEM_ADDR_WIDTH)
        port map (
            clk   => clk,
            wen   => op_addr_gen_wr_en,    -- TODO: connect to output address generator //DONE
            waddr => op_addr_gen_wr_addr,  -- TODO: connect to output address generator //DONE
            wdata => mux2_out(C_MEM_OUT_WIDTH-1 downto 0),  -- TODO: connect to pipeline output through mux //DONE
            raddr => mem_out_rd_addr,
            rdata => mem_out_rd_data);
	------------------------------------------------------------------------------
				
end default;
