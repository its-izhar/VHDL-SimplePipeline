-- Izhar Shaikh
-- File: controller.vhd
--
-- Description: Implements a Controller to control, which will in-turn control address generator, Block RAMs and pipeline. 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.config_pkg.all;
use work.user_pkg.all;

entity controller is

  port(clk      : in std_logic;
       rst      : in std_logic;
       
       -- Mode control out for address generators
       ip_addr_gen_mode_out 	: out std_logic;     -- 0: Read Mode, 1: Write Mode
	   op_addr_gen_mode_out		: out std_logic;
       
       -- Size of memory (i.e. The number of addressess to be generated by Address Generator)
       ip_addr_gen_size_out 	: out std_logic_vector(C_MEM_ADDR_WIDTH downto 0);
	   op_addr_gen_size_out 	: out std_logic_vector(C_MEM_ADDR_WIDTH downto 0);   
           
	   -- Address Generators Control I/O
       ip_addr_gen_go	    : out std_logic;
	   op_addr_gen_go	    : out std_logic;
       ip_addr_gen_done		: in std_logic;
	   op_addr_gen_done		: in std_logic;

       -- Controller Control I/O
       go    	: in std_logic;
       done  	: out std_logic;

	   -- Size in for controller
	   size		: in std_logic_vector(C_MEM_ADDR_WIDTH downto 0));   
	   
end controller;


architecture default of controller is
    
    type state_type is (S_WAIT_GO, S_INIT, S_INITIALIZE_ADDRESS_GENERATORS, S_START_ADDRESS_GENERATORS, S_WAIT_UNTIL_DONE, S_DONE);
    signal state : state_type;    
    
    constant C_READ_MODE : std_logic := '0';
    constant C_WRITE_MODE : std_logic := '1'; 
    
    signal regSize  : std_logic_vector(C_MEM_ADDR_WIDTH downto 0) := (others => '0');
    
begin
  process(clk, rst)
    
  begin

    if rst = '1' then
        state  <= S_WAIT_GO;
        done <= '0';
		-- Mode control out for address generators
		ip_addr_gen_mode_out <= C_READ_MODE;
		op_addr_gen_mode_out <= C_WRITE_MODE;     
		-- Size of memory (i.e. The number of addressess to be generated by Address Generator)
		ip_addr_gen_size_out <= (others => '0');
		op_addr_gen_size_out <= (others => '0');
		-- Address Generators Control I/O
		ip_addr_gen_go <= '0';
		op_addr_gen_go <= '0';
        
    elsif (rising_edge(clk)) then

        case state is
            when S_WAIT_GO =>
                if(go = '1') then
                    state <= S_INIT;
                end if;
                
            when S_INIT =>
				done <= '0';
				regSize <= size;
				state <= S_INITIALIZE_ADDRESS_GENERATORS;
				
			when S_INITIALIZE_ADDRESS_GENERATORS =>
				-- Mode control out for address generators
				ip_addr_gen_mode_out <= C_READ_MODE;
				op_addr_gen_mode_out <= C_WRITE_MODE;     
				-- Size of memory (i.e. The number of addressess to be generated by Address Generator)
				ip_addr_gen_size_out <= regSize;
				op_addr_gen_size_out <= regSize;
				-- Start the Addr Generators
				state <= S_START_ADDRESS_GENERATORS;
				
			when S_START_ADDRESS_GENERATORS =>
				-- Address Generators Control I/O
				ip_addr_gen_go <= '1';
				op_addr_gen_go <= '1';
                state <= S_WAIT_UNTIL_DONE;
                
            when S_WAIT_UNTIL_DONE =>
                if(ip_addr_gen_done = '1' and op_addr_gen_done = '1') then          -- Wait until both address generators are done
					done <= '1';
                    state <= S_DONE;
                end if;
                
            when S_DONE =>
                if (go = '0') then
                    state <= S_WAIT_GO;
                end if;
            
            when others =>
                NULL;
        
        end case;
    end if;
  end process; 
end default;
